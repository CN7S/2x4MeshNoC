module router_tb();
	







endmodule